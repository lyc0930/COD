`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/05/04 23:43:54
// Design Name: 
// Module Name: Hex7SegmentDisplay
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Hex7SegmentDisplay(x, seg);
    input  [3:0] x;
    output [6:0] seg; 
//                   0                                 1                                 2                                 3                                 4                                 5                                 6                                 7                                 8                                 9                                 A                                 b                                 C                                 d                                 E                                 F
//	assign AbCdEF = (~x[3] & ~x[2] & ~x[1] & ~x[0]) | (~x[3] & ~x[2] & ~x[1] &  x[0]) | (~x[3] & ~x[2] &  x[1] & ~x[0]) | (~x[3] & ~x[2] &  x[1] &  x[0]) | (~x[3] &  x[2] & ~x[1] & ~x[0]) | (~x[3] &  x[2] & ~x[1] &  x[0]) | (~x[3] &  x[2] &  x[1] & ~x[0]) | (~x[3] &  x[2] &  x[1] &  x[0]) | ( x[3] & ~x[2] & ~x[1] & ~x[0]) | ( x[3] & ~x[2] & ~x[1] &  x[0]) | ( x[3] & ~x[2] &  x[1] & ~x[0]) | ( x[3] & ~x[2] &  x[1] &  x[0]) | ( x[3] &  x[2] & ~x[1] & ~x[0]) | ( x[3] &  x[2] & ~x[1] &  x[0]) | ( x[3] &  x[2] &  x[1] & ~x[0]) | ( x[3] &  x[2] &  x[1] &  x[0]);
    assign seg[0] =                                   (~x[3] & ~x[2] & ~x[1] &  x[0]) |                                                                                                                                                                                                                                                                                                                   ( x[3] & ~x[2] &  x[1] &  x[0]) |                                   ( x[3] &  x[2] & ~x[1] &  x[0])                                                                    ;
    assign seg[1] =                                                                                                                                                                           (~x[3] &  x[2] & ~x[1] &  x[0]) | (~x[3] &  x[2] &  x[1] & ~x[0]) |                                                                                                                                         ( x[3] & ~x[2] &  x[1] &  x[0]) | ( x[3] &  x[2] & ~x[1] & ~x[0]) |                                   ( x[3] &  x[2] &  x[1] & ~x[0]) | ( x[3] &  x[2] &  x[1] &  x[0]);
    assign seg[2] =                                                                     (~x[3] & ~x[2] &  x[1] & ~x[0]) |                                                                                                                                                                                                                                                                                                                   ( x[3] &  x[2] & ~x[1] & ~x[0]) |                                   ( x[3] &  x[2] &  x[1] & ~x[0]) | ( x[3] &  x[2] &  x[1] &  x[0]);
    assign seg[3] =                                   (~x[3] & ~x[2] & ~x[1] &  x[0]) |                                                                     (~x[3] &  x[2] & ~x[1] & ~x[0]) |                                                                     (~x[3] &  x[2] &  x[1] &  x[0]) |                                   ( x[3] & ~x[2] & ~x[1] &  x[0]) | ( x[3] & ~x[2] &  x[1] & ~x[0]) |                                                                                                                                         ( x[3] &  x[2] &  x[1] &  x[0]);
    assign seg[4] =                                   (~x[3] & ~x[2] & ~x[1] &  x[0]) |                                   (~x[3] & ~x[2] &  x[1] &  x[0]) | (~x[3] &  x[2] & ~x[1] & ~x[0]) | (~x[3] &  x[2] & ~x[1] &  x[0]) |                                   (~x[3] &  x[2] &  x[1] &  x[0]) |                                   ( x[3] & ~x[2] & ~x[1] &  x[0])                                                                                                                                                                                                            ;
    assign seg[5] =                                   (~x[3] & ~x[2] & ~x[1] &  x[0]) | (~x[3] & ~x[2] &  x[1] & ~x[0]) | (~x[3] & ~x[2] &  x[1] &  x[0]) |                                                                                                       (~x[3] &  x[2] &  x[1] &  x[0]) |                                                                                                                                                                           ( x[3] &  x[2] & ~x[1] &  x[0])                                                                    ;
    assign seg[6] = (~x[3] & ~x[2] & ~x[1] & ~x[0]) | (~x[3] & ~x[2] & ~x[1] &  x[0]) |                                                                                                                                                                           (~x[3] &  x[2] &  x[1] &  x[0]) |                                                                                                                                         ( x[3] &  x[2] & ~x[1] & ~x[0])                                                                                                      ;  
endmodule

